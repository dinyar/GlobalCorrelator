library ieee;
use ieee.std_logic_1164.all;

package board_constants is
    constant N_QUADS : natural := 19;
end;
