library ieee;
use ieee.std_logic_1164.all;

package ultra_constants is
    constant N_QUADS : natural := 76;
end;

