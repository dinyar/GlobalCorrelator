library ieee;
use ieee.std_logic_1164.all;

package ultra_constants is
    constant DUMMY_ANSWER : natural := 42;
end;

